** Profile: "stab2Prot2-DC_Sweep_vI"  [ C:\Users\mvman\projects2\OrCAD\AnaSim\stabilizTensiune\stab_v1-stab2prot2-dc_sweep_vi.sim ] 

** Creating circuit file "stab_v1-stab2prot2-dc_sweep_vi.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 10 15 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\stab_v1-stab2Prot2.net" 


.END
