** Profile: "stab1RedrMono1-tran1"  [ C:\Users\mvman\projects2\OrCAD\AnaSim\stabilizTensiune\stab_v1-stab1RedrMono1-tran1.sim ] 

** Creating circuit file "stab_v1-stab1RedrMono1-tran1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.1s 0 1m 
.SAVEBIAS "C:\Users\mvman\projects2\OrCAD\AnaSim\stabilizTensiune\bias1" TRAN NOSUBCKT 
.OPTIONS LIST
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) 
.INC ".\stab_v1-stab1RedrMono1.net" 


.END
