** Profile: "stab1-DC_Sweep"  [ C:\Users\mvman\projects2\OrCAD\AnaSim\stabilizTensiune\stab_v1-stab1-dc_sweep.sim ] 

** Creating circuit file "stab_v1-stab1-dc_sweep.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 10 15 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\stab_v1-stab1.net" 


.END
